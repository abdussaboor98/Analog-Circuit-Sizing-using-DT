.param MOSFET_0_8_W_BIASCM_PMOS=4.2824265994131565 MOSFET_0_8_L_BIASCM_PMOS=1.774040549993515 MOSFET_0_8_M_BIASCM_PMOS=1
.param MOSFET_8_2_W_gm1_PMOS=6.452906936407089 MOSFET_8_2_L_gm1_PMOS=2.788204960525036 MOSFET_8_2_M_gm1_PMOS=9
.param MOSFET_10_1_W_gm2_PMOS=6.760543689131737 MOSFET_10_1_L_gm2_PMOS=3.273772805929184 MOSFET_10_1_M_gm2_PMOS=32
.param MOSFET_11_1_W_gmf2_PMOS=6.165277853608131 MOSFET_11_1_L_gmf2_PMOS=2.843104414641857 MOSFET_11_1_M_gmf2_PMOS=197
.param MOSFET_17_7_W_BIASCM_NMOS=8.30527549982071 MOSFET_17_7_L_BIASCM_NMOS=2.8800555169582367 MOSFET_17_7_M_BIASCM_NMOS=26
.param MOSFET_21_2_W_LOAD2_NMOS=3.877997562289238 MOSFET_21_2_L_LOAD2_NMOS=2.1998604550026357 MOSFET_21_2_M_LOAD2_NMOS=30
.param MOSFET_23_1_W_gm3_NMOS=3.782426029443741 MOSFET_23_1_L_gm3_NMOS=2.8648027116432786 MOSFET_23_1_M_gm3_NMOS=14
.param CURRENT_0_BIAS=1.679703786969185e-05
.param M_C0=42
.param M_C1=20
